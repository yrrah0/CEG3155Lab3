library verilog;
use verilog.vl_types.all;
entity testBench_vlg_vec_tst is
end testBench_vlg_vec_tst;
