library verilog;
use verilog.vl_types.all;
entity trafficlight_vlg_vec_tst is
end trafficlight_vlg_vec_tst;
